// List of RISC-V opcodes and funct codes.
// Use `include "Opcode.vh" to use these in the decoder

`ifndef OPCODE
`define OPCODE

// ***** Opcodes *****
// Special immediate instructions
`define OPC_LUI         7'b0110111
`define OPC_AUIPC       7'b0010111

// Jump instructions
`define OPC_JAL         7'b1101111
`define OPC_JALR        7'b1100111

// Branch instructions
`define OPC_BRANCH      7'b1100011

// Load and store instructions
`define OPC_STORE       7'b0100011
`define OPC_LOAD        7'b0000011

// Arithmetic instructions
`define OPC_ARI_RTYPE   7'b0110011
`define OPC_ARI_ITYPE   7'b0010011

// ***** 5-bit Opcodes *****
`define OPC_LUI_5       5'b01101
`define OPC_AUIPC_5     5'b00101
`define OPC_JAL_5       5'b11011
`define OPC_JALR_5      5'b11001
`define OPC_BRANCH_5    5'b11000
`define OPC_STORE_5     5'b01000
`define OPC_LOAD_5      5'b00000
`define OPC_ARI_RTYPE_5 5'b01100
`define OPC_ARI_ITYPE_5 5'b00100

// ***** Function codes *****

// Branch function codes
`define FNC_BEQ         3'b000
`define FNC_BNE         3'b001
`define FNC_BLT         3'b100
`define FNC_BGE         3'b101
`define FNC_BLTU        3'b110
`define FNC_BGEU        3'b111

// Load and store function codes
`define FNC_LB          3'b000
`define FNC_LH          3'b001
`define FNC_LW          3'b010
`define FNC_LBU         3'b100
`define FNC_LHU         3'b101
`define FNC_SB          3'b000
`define FNC_SH          3'b001
`define FNC_SW          3'b010

// Arithmetic R-type and I-type functions codes
`define FNC_ADD_SUB     3'b000
`define FNC_SLL         3'b001
`define FNC_SLT         3'b010
`define FNC_SLTU        3'b011
`define FNC_XOR         3'b100
`define FNC_OR          3'b110
`define FNC_AND         3'b111
`define FNC_SRL_SRA     3'b101

// ADD and SUB use the same opcode + function code
// SRA and SRL also use the same opcode + function code
// For these operations, we also need to look at bit 30 of the instruction
`define FNC2_ADD        1'b0
`define FNC2_SUB        1'b1
`define FNC2_SRL        1'b0
`define FNC2_SRA        1'b1

//my definition of opcode
`define LUI_OP 7'b0110111
`define AUIPC_OP 7'b0010111
`define JAL_OP 7'b1101111
`define JALR_OP 7'b1100111

`define BRANCH_OP 7'b1100011

`define LOARD_OP 7'b0000011

`define STORE_OP 7'b0100011

`define ARITH_IMM_OP 7'b0010011

`define ARITH_REG_OP 7'b0110011

`define CSR_OP 7'b1110011
`define CSRRWI_FUNCT 3'b101
`define CSRRW_FUNCT 3'b001

`define BEQ_FUNCT 3'b000
`define BNE_FUNCT 3'b001
`define BLT_FUNCT 3'b100
`define BGE_FUNCT 3'b101
`define BLTU_FUNCT 3'b110
`define BGEU_FUNCT 3'b111


`define LB_FUNCT 3'b000
`define LH_FUNCT 3'b001
`define LW_FUNCT 3'b010
`define LBU_FUNCT 3'b100
`define LHU_FUNCT 3'b101

`define SB_FUNCT 3'b000
`define SH_FUNCT 3'b001
`define SW_FUNCT 3'b010


`define ADDI_FUNCT 3'b000
`define SLTI_FUNCT 3'b010
`define SLTIU_FUNCT 3'b011
`define XORI_FUNCT 3'b100
`define ORI_FUNCT 3'b110
`define ANDI_FUNCT 3'b111
`define SLLI_FUNCT 3'b001
`define SRLI_FUNCT 3'b101
`define SRAI_FUNCT 3'b101

`define ADD_FUNCT 3'b000
`define SLL_FUNCT 3'b001
`define SLT_FUNCT 3'b010
`define SLTU_FUNCT 3'b011
`define XOR_FUNCT 3'b100
`define SRL_FUNCT 3'b101
`define OR_FUNCT 3'b110
`define AND_FUNCT 3'b111
`endif //OPCODE
